** Library name: ECE555
** Cell name: OR
** View name: schematic
mp4 y net2 vdd vdd pmos_lvt w=27e-9 l=20e-9 nfin=1
mp1 net2 b net1 net2 pmos_lvt w=27e-9 l=20e-9 nfin=1
mp0 net1 a vdd net2 pmos_lvt w=27e-9 l=20e-9 nfin=1
mn5 y net2 vss vss nmos_lvt w=27e-9 l=20e-9 nfin=1
mn3 net2 b vss vss nmos_lvt w=27e-9 l=20e-9 nfin=1
mn2 net2 a vss vss nmos_lvt w=27e-9 l=20e-9 nfin=1
.END
